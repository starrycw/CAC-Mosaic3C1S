`ifndef __TNS_HEADER__
    `define __TNS_HEADER__
    
    // TNS
    `define TNS01_C     1
    `define TNS01_B     2
    `define TNS01_A     3
    
    `define TNS02_C     7
    `define TNS02_B     14
    `define TNS02_A     21
    
    `define TNS03_C     49
    `define TNS03_B     98
    `define TNS03_A     147
    
    `define TNS04_C     343
    `define TNS04_B     686
    `define TNS04_A     1029
    
    `define TNS05_C     2401
    `define TNS05_B     4802
    `define TNS05_A     7203
    
    `define TNS06_C     16807
    `define TNS06_B     33614
    `define TNS06_A     50421
    
    `define TNS07_C     117649
    `define TNS07_B     235298
    `define TNS07_A     352947
    
    `define TNS08_C      823543
    `define TNS08_B      1647086
    `define TNS08_A      2470629
    
    `define TNS09_C      5764801
    `define TNS09_B      11529602
    `define TNS09_A      17294403
    
    `define TNS10_C      40353607
    `define TNS10_B      80707214
    `define TNS10_A      121060821
    
    `define TNS11_C      282475249
    `define TNS11_B      564950498
    `define TNS11_A      847425747

    `define TNS12_C      1977326743
    `define TNS12_B      3954653486
    `define TNS12_A      5931980229
    
    `define TNS13_C      13841287201
    `define TNS13_B      27682574402
    `define TNS13_A      41523861603
    
    `define TNS14_C      96889010407
    `define TNS14_B      193778020814
    `define TNS14_A      290667031221
    
    `define TNS15_C      678223072849
    `define TNS15_B      1356446145698
    `define TNS15_A      2034669218547
    
    `define TNS16_C      4747561509943
    `define TNS16_B      9495123019886
    `define TNS16_A      14242684529829


    

    //binary code len (eg: data[`BLEN_03-1 : 0] can be coded as 3-group TNS-CAC codewords)
    `define BLEN01_C    1
    `define BLEN01_B    2
    `define BLEN01      2
    
    `define BLEN02_C    3
    `define BLEN02_B    4
    `define BLEN02      5
    
    `define BLEN03_C    6
    `define BLEN03_B    7
    `define BLEN03      8
    
    `define BLEN04_C    9
    `define BLEN04_B    10
    `define BLEN04      11
    
    `define BLEN05_C    12
    `define BLEN05_B    13
    `define BLEN05      14
    
    `define BLEN06_C    15
    `define BLEN06_B    16
    `define BLEN06      16
    
    `define BLEN07_C    17
    `define BLEN07_B    18
    `define BLEN07      19
    
    `define BLEN08_C    20
    `define BLEN08_B    21
    `define BLEN08      22
    
    `define BLEN09_C    23
    `define BLEN09_B    24
    `define BLEN09      25
    
    `define BLEN10_C    26
    `define BLEN10_B    27
    `define BLEN10      28
    
    `define BLEN11_C    29
    `define BLEN11_B    30
    `define BLEN11      30
    
    `define BLEN12_C    31
    `define BLEN12_B    32
    `define BLEN12      33
    
    `define BLEN13_C    34
    `define BLEN13_B    35
    `define BLEN13      36
    
    `define BLEN14_C    37
    `define BLEN14_B    38
    `define BLEN14      39
    
    `define BLEN15_C    40
    `define BLEN15_B    41
    `define BLEN15      42
    
    `define BLEN16_C    43
    `define BLEN16_B    44
    `define BLEN16      44

    
    
    
    
    
    //remaining value len 
    `define RLEN01_C    1
    `define RLEN01_B    2
    `define RLEN01      3
    
    `define RLEN02_C    4
    `define RLEN02_B    5
    `define RLEN02      6
    
    `define RLEN03_C    7
    `define RLEN03_B    8
    `define RLEN03      9
    
    `define RLEN04_C    10
    `define RLEN04_B    11
    `define RLEN04      12
    
    `define RLEN05_C    13
    `define RLEN05_B    14
    `define RLEN05      15
    
    `define RLEN06_C    16
    `define RLEN06_B    17
    `define RLEN06      17
    
    `define RLEN07_C    18
    `define RLEN07_B    19
    `define RLEN07      20

    `define RLEN08_C    21
    `define RLEN08_B    22
    `define RLEN08      23
    
    `define RLEN09_C    24
    `define RLEN09_B    25
    `define RLEN09      26
    
    `define RLEN10_C    27
    `define RLEN10_B    28
    `define RLEN10      29
    
    `define RLEN11_C    30
    `define RLEN11_B    31
    `define RLEN11      31
    
    `define RLEN12_C    32
    `define RLEN12_B    33
    `define RLEN12      34
    
    `define RLEN13_C    35
    `define RLEN13_B    36
    `define RLEN13      37
    
    `define RLEN14_C    38
    `define RLEN14_B    39
    `define RLEN14      40
    
    `define RLEN15_C    41
    `define RLEN15_B    42
    `define RLEN15      43
    
    `define RLEN16_C    44
    `define RLEN16_B    45
    `define RLEN16      45

    
    
`endif
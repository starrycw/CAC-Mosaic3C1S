`ifndef __FNS_HEADER__
    `define __FNS_HEADER__
    
    //FNS
    `define FNS01   1
    `define FNS02   1
    `define FNS03   2
    `define FNS04   3
    `define FNS05   5
    `define FNS06   8
    `define FNS07   13
    `define FNS08   21
    `define FNS09   34
    `define FNS10   55
    `define FNS11   89
    `define FNS12   144
    `define FNS13   233
    `define FNS14   377
    `define FNS15   610
    `define FNS16   987
    `define FNS17   1597
    `define FNS18   2584
    `define FNS19   4181
    `define FNS20   6765
    `define FNS21   10946
    `define FNS22   17711
    `define FNS23   28657
    `define FNS24   46368
    `define FNS25   75025
    `define FNS26   121393
    `define FNS27   196418
    `define FNS28   317811
    `define FNS29   514229
    `define FNS30   832040
    `define FNS31   1346269
    `define FNS32   2178309
    `define FNS33   3524578
    `define FNS34   5702887
    `define FNS35   9227465
    `define FNS36   14930352
    `define FNS37   24157817
    `define FNS38   39088169
    `define FNS39   63245986
    `define FNS40   102334155
    `define FNS41   165580141
    `define FNS42   267914296
    `define FNS43   433494437
    `define FNS44   701408733
    `define FNS45   1134903170
    `define FNS46   1836311903



    `define FBLEN01  1
    `define FBLEN02  1
    `define FBLEN03  2
    `define FBLEN04  3
    `define FBLEN05  3
    `define FBLEN06  4
    `define FBLEN07  5
    `define FBLEN08  5
    `define FBLEN09  6
    `define FBLEN10  7
    `define FBLEN11  7
    `define FBLEN12  8
    `define FBLEN13  9
    `define FBLEN14  9
    `define FBLEN15  10
    `define FBLEN16  11
    `define FBLEN17  12
    `define FBLEN18  12
    `define FBLEN19  13
    `define FBLEN20  14
    `define FBLEN21  14
    `define FBLEN22  15
    `define FBLEN23  16
    `define FBLEN24  16
    `define FBLEN25  17
    `define FBLEN26  18
    `define FBLEN27  18
    `define FBLEN28  19
    `define FBLEN29  20   
    `define FBLEN30  21
    `define FBLEN31  21
    `define FBLEN32  22
    `define FBLEN33  23
    `define FBLEN34  23
    `define FBLEN35  24
    `define FBLEN36  25
    `define FBLEN37  25
    `define FBLEN38  26
    `define FBLEN39  27
    `define FBLEN40  27
    `define FBLEN41  28
    `define FBLEN42  29
    `define FBLEN43  30
    `define FBLEN44  30
    `define FBLEN45  31
    `define FBLEN46  32


    
    `define FRLEN01  1
    `define FRLEN02  2
    `define FRLEN03  3
    `define FRLEN04  3
    `define FRLEN05  4
    `define FRLEN06  5
    `define FRLEN07  6
    `define FRLEN08  6
    `define FRLEN09  7
    `define FRLEN10  8
    `define FRLEN11  8
    `define FRLEN12  9
    `define FRLEN13  10
    `define FRLEN14  10
    `define FRLEN15  11
    `define FRLEN16  12
    `define FRLEN17  13
    `define FRLEN18  13
    `define FRLEN19  14
    `define FRLEN20  15
    `define FRLEN21  15
    `define FRLEN22  16
    `define FRLEN23  17
    `define FRLEN24  17
    `define FRLEN25  18
    `define FRLEN26  19
    `define FRLEN27  19
    `define FRLEN28  20
    `define FRLEN29  21
    `define FRLEN30  22
    `define FRLEN31  22
    `define FRLEN32  23
    `define FRLEN33  24
    `define FRLEN34  24
    `define FRLEN35  25
    `define FRLEN36  26
    `define FRLEN37  26
    `define FRLEN38  27
    `define FRLEN39  28
    `define FRLEN40  28
    `define FRLEN41  29
    `define FRLEN42  30
    `define FRLEN43  31
    `define FRLEN44  31
    `define FRLEN45  32
    `define FRLEN46  33

    
    
    `define DBLEN01     1
    `define DBLEN02     2
    `define DBLEN03     2
    `define DBLEN04     3
    `define DBLEN05     4
    `define DBLEN06     4
    `define DBLEN07     5
    `define DBLEN08     6
    `define DBLEN09     6
    `define DBLEN10     7
    `define DBLEN11     8
    `define DBLEN12     8
    `define DBLEN13     9
    `define DBLEN14     10
    `define DBLEN15     10
    `define DBLEN16     11
    `define DBLEN17     12
    `define DBLEN18     13
    `define DBLEN19     13
    `define DBLEN20     14
    `define DBLEN21     15
    `define DBLEN22     15
    `define DBLEN23     16
    `define DBLEN24     17
    `define DBLEN25     17
    `define DBLEN26     18
    `define DBLEN27     19
    `define DBLEN28     19
    `define DBLEN29     20
    `define DBLEN30     21
    `define DBLEN31     22
    `define DBLEN32     22
    `define DBLEN33     23
    `define DBLEN34     24
    `define DBLEN35     24
    `define DBLEN36     25
    `define DBLEN37     26
    `define DBLEN38     26
    `define DBLEN39     27
    `define DBLEN40     28
    `define DBLEN41     28
    `define DBLEN42     29
    `define DBLEN43     30
    `define DBLEN44     31
    `define DBLEN45     31
    `define DBLEN46     32


    `define DRLEN01     1
    `define DRLEN02     2
    `define DRLEN03     3
    `define DRLEN04     4
    `define DRLEN05     4
    `define DRLEN06     5
    `define DRLEN07     6
    `define DRLEN08     7
    `define DRLEN09     7
    `define DRLEN10     8
    `define DRLEN11     9
    `define DRLEN12     9
    `define DRLEN13     10
    `define DRLEN14     11
    `define DRLEN15     11
    `define DRLEN16     12
    `define DRLEN17     13
    `define DRLEN18     14
    `define DRLEN19     14
    `define DRLEN20     15
    `define DRLEN21     16
    `define DRLEN22     16
    `define DRLEN23     17
    `define DRLEN24     18
    `define DRLEN25     18
    `define DRLEN26     19
    `define DRLEN27     20
    `define DRLEN28     20
    `define DRLEN29     21
    `define DRLEN30     22
    `define DRLEN31     23
    `define DRLEN32     23
    `define DRLEN33     24
    `define DRLEN34     25
    `define DRLEN35     25
    `define DRLEN36     26
    `define DRLEN37     27
    `define DRLEN38     27
    `define DRLEN39     28
    `define DRLEN40     29
    `define DRLEN41     29
    `define DRLEN42     30
    `define DRLEN43     31
    `define DRLEN44     32
    `define DRLEN45     32
    `define DRLEN46     33

    
    `define IBLEN01     1
    `define IBLEN02     1
    `define IBLEN03     2
    `define IBLEN04     3
    `define IBLEN05     4
    `define IBLEN06     4
    `define IBLEN07     5
    `define IBLEN08     6
    `define IBLEN09     6
    `define IBLEN10     7
    `define IBLEN11     8
    `define IBLEN12     8
    `define IBLEN13     9
    `define IBLEN14     10
    `define IBLEN15     10
    `define IBLEN16     11
    `define IBLEN17     12
    `define IBLEN18     13
    `define IBLEN19     13
    `define IBLEN20     14
    `define IBLEN21     15
    `define IBLEN22     15
    `define IBLEN23     16
    `define IBLEN24     17
    `define IBLEN25     17
    `define IBLEN26     18
    `define IBLEN27     19
    `define IBLEN28     19
    `define IBLEN29     20
    `define IBLEN30     21
    `define IBLEN31     22
    `define IBLEN32     22
    `define IBLEN33     23
    `define IBLEN34     24
    `define IBLEN35     24
    `define IBLEN36     25
    `define IBLEN37     26
    `define IBLEN38     26
    `define IBLEN39     27
    `define IBLEN40     28
    `define IBLEN41     28
    `define IBLEN42     29
    `define IBLEN43     30
    `define IBLEN44     31
    `define IBLEN45     31
    `define IBLEN46     32

    
    
    `define IRLEN01     1
    `define IRLEN02     2
    `define IRLEN03     3
    `define IRLEN04     4
    `define IRLEN05     4
    `define IRLEN06     5
    `define IRLEN07     6
    `define IRLEN08     7
    `define IRLEN09     7
    `define IRLEN10     8
    `define IRLEN11     9
    `define IRLEN12     9
    `define IRLEN13     10
    `define IRLEN14     11
    `define IRLEN15     11
    `define IRLEN16     12
    `define IRLEN17     13
    `define IRLEN18     14
    `define IRLEN19     14
    `define IRLEN20     15
    `define IRLEN21     16
    `define IRLEN22     16
    `define IRLEN23     17
    `define IRLEN24     18
    `define IRLEN25     18
    `define IRLEN26     19
    `define IRLEN27     20
    `define IRLEN28     20
    `define IRLEN29     21
    `define IRLEN30     22
    `define IRLEN31     23
    `define IRLEN32     23
    `define IRLEN33     24
    `define IRLEN34     25
    `define IRLEN35     25
    `define IRLEN36     26
    `define IRLEN37     27
    `define IRLEN38     27
    `define IRLEN39     28
    `define IRLEN40     29
    `define IRLEN41     29
    `define IRLEN42     30
    `define IRLEN43     31
    `define IRLEN44     32
    `define IRLEN45     32
    `define IRLEN46     33








    
    
    
`endif
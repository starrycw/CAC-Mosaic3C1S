//  ������ϵCAC����
//  
//  1. Design Sources
//  
//      1.1 TNS.vh
//          ��TNS��ϵ�йصĶ���
//      1.2 FNS.vh
//          ��FNS��ϵ�йصĶ��壬�Լ���IDP/3D-DPS�����йصĶ���
//      1.3 TNS_encoder_xx/TNS_dec_xx
//          TNS���������xxΪ���볤��
//      1.4 FPF_encoder_xx/FNS_dec_xx
//          FNS FPF���������xxΪ���볤��
//      1.5 FTF_encoder_xx/FNS_dec_xx
//          FNS FTF���������xxΪ���볤��
//      1.6 IDP_encoder_xx/IDP_dec_xx
//          IDP���������xxΪ���볤��
//      1.7 DPS_encoder_xx/DPS_dec_xx
//          3D-DPS���������xxΪ���볤��
//  2. Simulation Sources
//
//      2.1 Simu_TNS_xx
//          ��֤TNS����빦��
//      2.2 Simu_FPF_xx
//          ��֤FPF����빦��
//      2.3 Simu_FTF_xx
//          ��֤FTF����빦��
//      2.4 Simu_IDP_xx
//          ��֤IDP����빦��
//      2.5 Simu_DPS_xx
//          ��֤3D-DPS����빦��
//
//
//
//  3. Revision
//
//      ��2020.05.14�� - ����
//      ��2020.06.06�� - ���벿�ֳ��ȵ�����ʱ�����ֱ����������С���ֳ���
//                          Datalen:    5   8   11  14  17  20  23  26  29
//                          TNS:        6   9   12  15  19  22  25  28  31
//                          FNS:        7   12  16  20  25  29  33  38  42
//                          3DDPS:      7   11  16  20  24  29  33  37  42
//                          IDP:        7   11  16  20  24  29  33  37  42